module core_top
(
    input           aclk,
    input           aresetn,
    input    [ 7:0] intrpt, 
    output   [ 3:0] arid,
    output   [31:0] araddr,
    output   [ 7:0] arlen,
    output   [ 2:0] arsize,
    output   [ 1:0] arburst,
    output   [ 1:0] arlock,
    output   [ 3:0] arcache,
    output   [ 2:0] arprot,
    output          arvalid,
    input           arready,
    input    [ 3:0] rid,
    input    [31:0] rdata,
    input    [ 1:0] rresp,
    input           rlast,
    input           rvalid,
    output          rready,
    output   [ 3:0] awid,
    output   [31:0] awaddr,
    output   [ 7:0] awlen,
    output   [ 2:0] awsize,
    output   [ 1:0] awburst,
    output   [ 1:0] awlock,
    output   [ 3:0] awcache,
    output   [ 2:0] awprot,
    output          awvalid,
    input           awready,
    output   [ 3:0] wid,
    output   [31:0] wdata,
    output   [ 3:0] wstrb,
    output          wlast,
    output          wvalid,
    input           wready,
    input    [ 3:0] bid,
    input    [ 1:0] bresp,
    input           bvalid,
    output          bready
);

mycpu_top inner_cpu(
  .aclk(aclk),
  .aresetn(aresetn),
  .ext_int(intrpt),
  .awvalid(awvalid),
  .awready(awready),
  .awaddr(awaddr),
  .awid(awid),
  .awlen(awlen),
  .awsize(awsize),
  .awburst(awburst),
  .awlock(awlock),
  .awcache(awcache),
  .awprot(awprot),
  .wvalid(wvalid),
  .wready(wready),
  .wdata(wdata),
  .wstrb(wstrb),
  .wlast(wlast),
  .bvalid(bvalid),
  .bready(bready),
  .bid(bid),
  .bresp(bresp),
  .arvalid(arvalid),
  .arready(arready),
  .araddr(araddr),
  .arid(arid),
  .arlen(arlen),
  .arsize(arsize),
  .arburst(arburst),
  .arlock(arlock),
  .arcache(arcache),
  .arprot(arprot),
  .rvalid(rvalid),
  .rready(rready),
  .rdata(rdata),
  .rid(rid),
  .rresp(rresp),
  .rlast(rlast),
  .wid(wid)
);

endmodule